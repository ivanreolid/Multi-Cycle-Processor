`include "config.svh"

package params_pkg;

  parameter int OPCODE_WIDTH     = 4;
  parameter int REGISTER_WIDTH   = 5;
  parameter int SHAMT_WIDTH      = 6;
  parameter int CSR_ADDR_WIDTH   = 12;
  parameter int INSTR_WIDTH      = 32;
  parameter int ADDR_WIDTH       = 32;
  parameter int DATA_WIDTH       = 32;
  parameter int MEM_SIZE         = 200000;

  parameter int ROB_ENTRIES      = `ROB_ENTRIES_MACRO;
  parameter int ROB_ENTRY_WIDTH  = $clog2(ROB_ENTRIES);

  parameter int VADDR_WIDTH       = 32;
  parameter int PADDR_WIDTH       = 20;
  parameter int PAGE_OFFSET_WIDTH = 12;
  parameter int VPN_WIDTH         = VADDR_WIDTH - PAGE_OFFSET_WIDTH;
  parameter int PPN_WIDTH         = PADDR_WIDTH - PAGE_OFFSET_WIDTH;

  parameter int ITLB_DEPTH       = `ITLB_DEPTH_MACRO;

  parameter int CACHE_LINE_BYTES = `CACHE_LINE_BYTES_MACRO;
  parameter int DCACHE_N_LINES   = `DCACHE_N_LINES_MACRO;
  parameter int ICACHE_N_LINES   = `ICACHE_N_LINES_MACRO;

  // CSRS
  parameter int CSR_SATP = 12'h180;

  typedef enum logic[6:0] {
    R         = 7'b0110011,
    LOAD      = 7'b0000011,
    STORE     = 7'b0100011,
    BRANCH    = 7'b1100011,
    JAL       = 7'b1101111,
    IMMEDIATE = 7'b0010011,
    LUI       = 7'b0110111,
    AUIPC     = 7'b0010111,
    SYSTEM    = 7'b1110011
  } opcode;

  typedef enum logic [2:0] {
    CSRRW = 3'b001
  } csr_op_t;

  typedef struct packed {
    logic is_mul;
    logic rs1_needed;
    logic rs2_needed;
    logic [4:0] rs1;
    logic [4:0] rs2;
  } hazard_ctrl_t;

  typedef enum logic [1:0] {
    BYTE  = 2'b00,
    HALF  = 2'b01,
    WORD  = 2'b10
  } access_size_t;

  function string opcode_to_string(opcode op);
    case (op)
      R         : opcode_to_string = "R";
      LOAD      : opcode_to_string = "LOAD";
      STORE     : opcode_to_string = "STORE";
      BRANCH    : opcode_to_string = "BRANCH";
      JAL       : opcode_to_string = "JAL";
      IMMEDIATE : opcode_to_string = "IMMEDIATE";
      LUI       : opcode_to_string = "LUI";
      AUIPC     : opcode_to_string = "AUIPC";
      SYSTEM    : opcode_to_string = "SYSTEM";
      default   : opcode_to_string = "???";
    endcase
  endfunction

  typedef struct packed {
    logic [6:0] funct7;
    logic [4:0] rs2;
    logic [4:0] rs1;
    logic [2:0] funct3;
    logic [4:0] rd;
    opcode opcode;
  } instruction_t;

endpackage
