`include "imem.sv"

import params_pkg::*;

module fetch_stage #(
  parameter int ADDR_WIDTH = params_pkg::ADDR_WIDTH,
  parameter int DATA_WIDTH = params_pkg::DATA_WIDTH,
  parameter int MEM_SIZE   = params_pkg::MEM_SIZE
)(
  input  logic clk_i,
  input  logic rst_i,
  input  logic alu_branch_taken_i,
  input  logic is_jump_i,
  input  logic [ADDR_WIDTH-1:0] pc_branch_offset_i,
  input  logic [ADDR_WIDTH-1:0] jump_address_i,
  input  logic instr_valid_i,
  input  instruction_t instr_i,
  output logic imem_req_valid_o,
  output logic dec_valid_o,
  output logic [ADDR_WIDTH-1:0] imem_req_pc_o,
  output logic [ADDR_WIDTH-1:0] dec_pc_o,
  output instruction_t instruction_o
);

  typedef enum logic [1:0] {
    IDLE     = 2'b00,
    MEM_REQ  = 2'b01,
    MEM_WAIT = 2'b10,
    FLUSH    = 2'b11
  } state_t;

  logic [ADDR_WIDTH-1:0] pc, pc_d, dec_pc_d;
  logic [ADDR_WIDTH-1:0] branch_target;

  state_t state, state_d;

  logic dec_valid_d;

  instruction_t dec_instr_d;

  always_comb begin : state_update
    imem_req_valid_o = 1'b0;
    imem_req_pc_o    = pc;
    dec_valid_d      = 1'b0;
    state_d          = state;
    pc_d             = pc;

    case (state)
      IDLE: begin
        state_d = MEM_REQ;
      end
      MEM_REQ: begin
        imem_req_valid_o = 1'b1;
        imem_req_pc_o    = pc;
        state_d          = MEM_WAIT;
      end
      MEM_WAIT: begin
        if (alu_branch_taken_i | is_jump_i)
          state_d = FLUSH;
        else if (instr_valid_i) begin
          dec_valid_d   = 1'b1;
          dec_instr_d   = instr_i;
          dec_pc_d      = pc;
          pc_d          = (pc + 1) % MEM_SIZE;
          state_d       = MEM_REQ;
        end
      end
      FLUSH: begin
        if (instr_valid_i) begin
          pc_d    = branch_target;
          state_d = MEM_REQ;
        end
      end
    endcase
  end

  always_ff @(posedge clk_i) begin : flops
    if (!rst_i) begin
      state          <= IDLE;
      pc             <= 1;
      branch_target  <= '0;
      dec_valid_o    <= 1'b0;
      dec_pc_o       <= '0;
      instruction_o  <= '0;
    end else begin
      state          <= state_d;
      pc             <= pc_d;
      dec_valid_o    <= dec_valid_d;
      dec_pc_o       <= dec_pc_d;
      instruction_o  <= dec_instr_d;

      if (alu_branch_taken_i)
        branch_target <= pc_branch_offset_i;
      else if (is_jump_i)
        branch_target <= jump_address_i;
    end
  end

endmodule : fetch_stage
